//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "FA4.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] w20;    //: /sn:0 {0}(#:658,268)(760,268)(#:760,194){1}
reg [3:0] w5;    //: /sn:0 {0}(#:367,111)(#:367,38){1}
wire [7:0] w7;    //: /sn:0 {0}(#:362,440)(362,478)(578,478)(578,424){1}
wire w14;    //: /sn:0 {0}(337,434)(337,417)(274,417)(274,351){1}
wire w16;    //: /sn:0 {0}(357,434)(357,383)(344,383)(344,351){1}
wire w15;    //: /sn:0 {0}(327,434)(327,423)(238,423)(238,351){1}
wire w4;    //: /sn:0 {0}(362,117)(362,149)(324,149)(324,172){1}
wire w19;    //: /sn:0 {0}(387,434)(387,417)(459,417)(459,351){1}
wire w0;    //: /sn:0 {0}(382,117)(382,134)(487,134)(487,172){1}
wire w3;    //: /sn:0 {0}(248,172)(248,132)(352,132)(352,117){1}
wire w1;    //: /sn:0 {0}(372,117)(372,149)(411,149)(411,172){1}
wire w8;    //: /sn:0 {0}(397,434)(397,423)(496,423)(496,351){1}
wire w30;    //: /sn:0 {0}(544,211)(637,211)(637,253)(652,253){1}
wire w17;    //: /sn:0 {0}(367,434)(367,383)(379,383)(379,351){1}
wire w10;    //: /sn:0 {0}(377,434)(377,409)(417,409)(417,351){1}
wire w13;    //: /sn:0 {0}(347,434)(347,409)(309,409)(309,351){1}
wire w27;    //: /sn:0 {0}(544,283)(597,283)(597,273)(652,273){1}
wire w29;    //: /sn:0 {0}(544,251)(596,251)(596,263)(652,263){1}
wire w26;    //: /sn:0 {0}(544,313)(637,313)(637,283)(652,283){1}
//: enddecls

  //: LED g4 (w7) @(578,417) /sn:0 /w:[ 1 ] /type:3
  //: DIP g3 (w20) @(760,184) /sn:0 /w:[ 1 ] /st:1 /dn:1
  assign {w30, w29, w27, w26} = w20; //: CONCAT g2  @(657,268) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  assign w7 = {w8, w19, w10, w17, w16, w13, w14, w15}; //: CONCAT g1  @(362,439) /sn:0 /R:3 /w:[ 0 0 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:1
  //: DIP g9 (w5) @(367,28) /sn:0 /w:[ 1 ] /st:2 /dn:1
  assign {w3, w4, w1, w0} = w5; //: CONCAT g17  @(367,112) /sn:0 /R:1 /w:[ 1 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  MUL g0 (.A3(w3), .A2(w4), .A1(w1), .A0(w0), .B0(w26), .B1(w27), .B2(w29), .B3(w30), .S0(w15), .S1(w14), .S2(w13), .S3(w16), .S4(w17), .S5(w10), .S6(w19), .S7(w8));   //: @(198, 173) /sz:(345, 177) /sn:0 /p:[ Ti0>0 Ti1>1 Ti2>1 Ti3>1 Ri0>0 Ri1>0 Ri2>0 Ri3>0 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<1 Bo6<1 Bo7<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FAb
module FAb(Cout, Cin, B, A, S);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(156,149)(201,149){1}
//: {2}(205,149)(227,149)(227,132)(242,132){3}
//: {4}(203,151)(203,281)(242,281){5}
input A;    //: /sn:0 {0}(156,118)(175,118){1}
//: {2}(179,118)(227,118)(227,127)(242,127){3}
//: {4}(177,120)(177,286)(242,286){5}
output Cout;    //: /sn:0 {0}(430,282)(511,282){1}
input Cin;    //: /sn:0 {0}(156,208)(251,208){1}
//: {2}(255,208)(394,208)(394,168)(409,168){3}
//: {4}(253,210)(253,241)(337,241){5}
output S;    //: /sn:0 {0}(430,166)(503,166){1}
wire w3;    //: /sn:0 {0}(358,239)(387,239)(387,279)(409,279){1}
wire w2;    //: /sn:0 {0}(263,130)(322,130)(322,161){1}
//: {2}(324,163)(367,163)(367,163)(409,163){3}
//: {4}(322,165)(322,236)(337,236){5}
wire w5;    //: /sn:0 {0}(263,284)(336,284)(336,284)(409,284){1}
//: enddecls

  _GGNAND2 #(4) g8 (.I0(w3), .I1(w5), .Z(Cout));   //: @(420,282) /sn:0 /w:[ 1 1 0 ]
  _GGNAND2 #(4) g4 (.I0(B), .I1(A), .Z(w5));   //: @(253,284) /sn:0 /w:[ 5 5 0 ]
  //: OUT g13 (Cout) @(508,282) /sn:0 /w:[ 1 ]
  _GGXOR2 #(8) g3 (.I0(A), .I1(B), .Z(w2));   //: @(253,130) /sn:0 /w:[ 3 3 0 ]
  //: IN g2 (Cin) @(154,208) /sn:0 /w:[ 0 ]
  //: IN g1 (B) @(154,149) /sn:0 /w:[ 0 ]
  //: joint g11 (Cin) @(253, 208) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g10 (.I0(w2), .I1(Cin), .Z(S));   //: @(420,166) /sn:0 /w:[ 3 3 0 ]
  //: joint g6 (B) @(203, 149) /w:[ 2 -1 1 4 ]
  //: joint g9 (w2) @(322, 163) /w:[ 2 1 -1 4 ]
  _GGNAND2 #(4) g7 (.I0(w2), .I1(Cin), .Z(w3));   //: @(348,239) /sn:0 /w:[ 5 5 0 ]
  //: joint g5 (A) @(177, 118) /w:[ 2 -1 1 4 ]
  //: IN g0 (A) @(154,118) /sn:0 /w:[ 0 ]
  //: OUT g12 (S) @(500,166) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FAdA
module FAdA(in4, C2, C1, in3);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output C2;    //: /sn:0 {0}(371,217)(260,217){1}
input in4;    //: /sn:0 {0}(134,142)(183,142){1}
//: {2}(187,142)(224,142)(224,114)(239,114){3}
//: {4}(185,144)(185,214)(239,214){5}
input in3;    //: /sn:0 {0}(134,85)(151,85){1}
//: {2}(155,85)(224,85)(224,109)(239,109){3}
//: {4}(153,87)(153,219)(239,219){5}
output C1;    //: /sn:0 {0}(260,112)(370,112){1}
//: enddecls

  //: joint g4 (in3) @(153, 85) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g3 (.I0(in4), .I1(in3), .Z(C2));   //: @(250,217) /sn:0 /w:[ 5 5 1 ]
  _GGXOR2 #(8) g2 (.I0(in3), .I1(in4), .Z(C1));   //: @(250,112) /sn:0 /w:[ 3 3 0 ]
  //: IN g1 (in4) @(132,142) /sn:0 /w:[ 0 ]
  //: OUT g6 (C2) @(368,217) /sn:0 /w:[ 0 ]
  //: OUT g7 (C1) @(367,112) /sn:0 /w:[ 1 ]
  //: joint g5 (in4) @(185, 142) /w:[ 2 -1 1 4 ]
  //: IN g0 (in3) @(132,85) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA3alt
module FA3alt(C1, Cin, C, B, S, C2, A);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(468,36)(526,36)(526,114){1}
input A;    //: /sn:0 {0}(418,68)(464,68)(464,114){1}
output C2;    //: /sn:0 {0}(121,349)(219,349){1}
input C;    //: /sn:0 {0}(469,307)(469,252)(425,252){1}
input Cin;    //: /sn:0 {0}(664,170)(560,170){1}
output C1;    //: /sn:0 {0}(283,455)(283,394){1}
output S;    //: /sn:0 {0}(503,452)(503,391){1}
wire w0;    //: /sn:0 {0}(517,307)(517,266)(501,266)(501,226){1}
wire w3;    //: /sn:0 {0}(442,349)(384,349)(384,264)(306,264)(306,307){1}
wire w1;    //: /sn:0 {0}(436,170)(248,170)(248,307){1}
//: enddecls

  FA g4 (.B(B), .A(A), .Cin(Cin), .Cout(w1), .Sin(w0));   //: @(437, 115) /sz:(122, 110) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: OUT g8 (C1) @(283,452) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (Cin) @(666,170) /sn:0 /R:2 /w:[ 0 ]
  //: IN g2 (C) @(423,252) /sn:0 /w:[ 1 ]
  //: IN g1 (B) @(466,36) /sn:0 /w:[ 0 ]
  //: OUT g6 (S) @(503,449) /sn:0 /R:3 /w:[ 0 ]
  FAdA g7 (.in4(w3), .in3(w1), .C2(C2), .C1(C1));   //: @(220, 308) /sz:(120, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: OUT g9 (C2) @(124,349) /sn:0 /R:2 /w:[ 0 ]
  FAd g5 (.in1(C), .in2(w0), .CoutFAd(w3), .S(S));   //: @(443, 308) /sz:(113, 82) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<1 ]
  //: IN g0 (A) @(416,68) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FAd
module FAd(in2, CoutFAd, S, in1);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(134,85)(151,85){1}
//: {2}(155,85)(224,85)(224,109)(239,109){3}
//: {4}(153,87)(153,219)(239,219){5}
input in2;    //: /sn:0 {0}(134,142)(183,142){1}
//: {2}(187,142)(224,142)(224,114)(239,114){3}
//: {4}(185,144)(185,214)(239,214){5}
output CoutFAd;    //: /sn:0 {0}(371,217)(260,217){1}
output S;    //: /sn:0 {0}(260,112)(370,112){1}
//: enddecls

  //: joint g4 (in1) @(153, 85) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g3 (.I0(in2), .I1(in1), .Z(CoutFAd));   //: @(250,217) /sn:0 /w:[ 5 5 1 ]
  _GGXOR2 #(8) g2 (.I0(in1), .I1(in2), .Z(S));   //: @(250,112) /sn:0 /w:[ 3 3 0 ]
  //: IN g1 (in2) @(132,142) /sn:0 /w:[ 0 ]
  //: OUT g6 (CoutFAd) @(368,217) /sn:0 /w:[ 0 ]
  //: OUT g7 (S) @(367,112) /sn:0 /w:[ 1 ]
  //: joint g5 (in2) @(185, 142) /w:[ 2 -1 1 4 ]
  //: IN g0 (in1) @(132,85) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA3b
module FA3b(C1, Cin, C, B, S, C2, A);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(468,36)(526,36)(526,114){1}
input A;    //: /sn:0 {0}(418,68)(464,68)(464,114){1}
output C2;    //: /sn:0 {0}(121,349)(219,349){1}
input C;    //: /sn:0 {0}(469,307)(469,252)(425,252){1}
input Cin;    //: /sn:0 {0}(664,170)(560,170){1}
output C1;    //: /sn:0 {0}(283,455)(283,394){1}
output S;    //: /sn:0 {0}(503,452)(503,391){1}
wire w0;    //: /sn:0 {0}(517,307)(517,266)(501,266)(501,226){1}
wire w3;    //: /sn:0 {0}(442,349)(384,349)(384,264)(306,264)(306,307){1}
wire w1;    //: /sn:0 {0}(436,170)(248,170)(248,307){1}
//: enddecls

  FA g4 (.B(B), .A(A), .Cin(Cin), .Cout(w1), .Sin(w0));   //: @(437, 115) /sz:(122, 110) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: OUT g8 (C1) @(283,452) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (Cin) @(666,170) /sn:0 /R:2 /w:[ 0 ]
  //: IN g2 (C) @(423,252) /sn:0 /w:[ 1 ]
  //: IN g1 (B) @(466,36) /sn:0 /w:[ 0 ]
  //: OUT g6 (S) @(503,449) /sn:0 /R:3 /w:[ 0 ]
  FAdA g7 (.in4(w3), .in3(w1), .C2(C2), .C1(C1));   //: @(220, 308) /sz:(120, 85) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: OUT g9 (C2) @(124,349) /sn:0 /R:2 /w:[ 0 ]
  FAd g5 (.in1(C), .in2(w0), .CoutFAd(w3), .S(S));   //: @(443, 308) /sz:(113, 82) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<1 ]
  //: IN g0 (A) @(416,68) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FAdD
module FAdD(in2, CoutFAd, S, in1);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(134,85)(151,85){1}
//: {2}(155,85)(224,85)(224,109)(239,109){3}
//: {4}(153,87)(153,219)(239,219){5}
input in2;    //: /sn:0 {0}(134,142)(183,142){1}
//: {2}(187,142)(224,142)(224,114)(239,114){3}
//: {4}(185,144)(185,214)(239,214){5}
output CoutFAd;    //: /sn:0 {0}(371,217)(260,217){1}
output S;    //: /sn:0 {0}(260,112)(370,112){1}
//: enddecls

  //: joint g4 (in1) @(153, 85) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g3 (.I0(in2), .I1(in1), .Z(CoutFAd));   //: @(250,217) /sn:0 /w:[ 5 5 1 ]
  _GGXOR2 #(8) g2 (.I0(in1), .I1(in2), .Z(S));   //: @(250,112) /sn:0 /w:[ 3 3 0 ]
  //: IN g1 (in2) @(132,142) /sn:0 /w:[ 0 ]
  //: OUT g6 (CoutFAd) @(368,217) /sn:0 /w:[ 0 ]
  //: OUT g7 (S) @(367,112) /sn:0 /w:[ 1 ]
  //: joint g5 (in2) @(185, 142) /w:[ 2 -1 1 4 ]
  //: IN g0 (in1) @(132,85) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUL
module MUL(S7, S2, S3, B3, B1, S1, B2, S4, S6, A0, A3, S0, A2, B0, A1, S5);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input A0;    //: /sn:0 {0}(-619,-207)(-353,-207){1}
//: {2}(-349,-207)(-6,-207){3}
//: {4}(-2,-207)(341,-207){5}
//: {6}(345,-207)(697,-207){7}
//: {8}(701,-207)(750,-207){9}
//: {10}(699,-205)(699,88){11}
//: {12}(343,-205)(343,55){13}
//: {14}(-4,-205)(-4,23){15}
//: {16}(-351,-205)(-351,-6){17}
output S1;    //: /sn:0 {0}(600,403)(600,462){1}
output S7;    //: /sn:0 {0}(-594,362)(-611,362)(-611,459){1}
output S6;    //: /sn:0 {0}(-452,408)(-452,433)(-452,433)(-452,459){1}
input A3;    //: /sn:0 {0}(-228,23)(-228,-84)(-228,-84)(-228,-97){1}
//: {2}(-226,-99)(117,-99){3}
//: {4}(121,-99)(473,-99){5}
//: {6}(477,-99)(753,-99){7}
//: {8}(475,-97)(475,88){9}
//: {10}(119,-97)(119,55){11}
//: {12}(-230,-99)(-573,-99){13}
//: {14}(-577,-99)(-619,-99){15}
//: {16}(-575,-97)(-575,-6){17}
input A2;    //: /sn:0 {0}(-619,-140)(-498,-140){1}
//: {2}(-494,-140)(-151,-140){3}
//: {4}(-147,-140)(196,-140){5}
//: {6}(200,-140)(552,-140){7}
//: {8}(556,-140)(751,-140){9}
//: {10}(554,-138)(554,88){11}
//: {12}(198,-138)(198,55){13}
//: {14}(-149,-138)(-149,23){15}
//: {16}(-496,-138)(-496,-6){17}
output S4;    //: /sn:0 {0}(-49,408)(-49,460){1}
input B2;    //: /sn:0 {0}(-263,-17)(-225,-17){1}
//: {2}(-221,-17)(-146,-17){3}
//: {4}(-142,-17)(-75,-17){5}
//: {6}(-71,-17)(-1,-17){7}
//: {8}(3,-17)(57,-17){9}
//: {10}(1,-15)(1,23){11}
//: {12}(-73,-15)(-73,23){13}
//: {14}(-144,-15)(-144,23){15}
//: {16}(-223,-15)(-223,23){17}
input B1;    //: /sn:0 {0}(84,15)(122,15){1}
//: {2}(126,15)(201,15){3}
//: {4}(205,15)(272,15){5}
//: {6}(276,15)(346,15){7}
//: {8}(350,15)(412,15){9}
//: {10}(348,17)(348,55){11}
//: {12}(274,17)(274,55){13}
//: {14}(203,17)(203,55){15}
//: {16}(124,17)(124,55){17}
output S0;    //: /sn:0 {0}(701,109)(701,459)(701,459)(701,462){1}
output S5;    //: /sn:0 {0}(-265,407)(-265,432)(-265,432)(-265,459){1}
input A1;    //: /sn:0 {0}(-620,-175)(-427,-175){1}
//: {2}(-423,-175)(-80,-175){3}
//: {4}(-76,-175)(267,-175){5}
//: {6}(271,-175)(623,-175){7}
//: {8}(627,-175)(750,-175){9}
//: {10}(625,-173)(625,88){11}
//: {12}(269,-173)(269,55){13}
//: {14}(-78,-173)(-78,23){15}
//: {16}(-425,-173)(-425,-6){17}
input B3;    //: /sn:0 {0}(-617,-46)(-572,-46){1}
//: {2}(-568,-46)(-493,-46){3}
//: {4}(-489,-46)(-422,-46){5}
//: {6}(-418,-46)(-348,-46){7}
//: {8}(-344,-46)(-297,-46){9}
//: {10}(-346,-44)(-346,-6){11}
//: {12}(-420,-44)(-420,-6){13}
//: {14}(-491,-44)(-491,-6){15}
//: {16}(-570,-44)(-570,-6){17}
output S3;    //: /sn:0 {0}(178,407)(178,462){1}
input B0;    //: /sn:0 {0}(439,49)(478,49){1}
//: {2}(482,49)(557,49){3}
//: {4}(561,49)(628,49){5}
//: {6}(632,49)(702,49){7}
//: {8}(706,49)(761,49){9}
//: {10}(704,51)(704,88){11}
//: {12}(630,51)(630,88){13}
//: {14}(559,51)(559,88){15}
//: {16}(480,51)(480,88){17}
output S2;    //: /sn:0 {0}(391,406)(391,462){1}
wire w32;    //: /sn:0 {0}(-226,44)(-226,81)(-266,81)(-266,307){1}
wire w6;    //: /sn:0 {0}(121,76)(121,112)(-29,112)(-29,293){1}
wire w7;    //: /sn:0 {0}(334,377)(293,377)(293,369)(248,369){1}
wire w16;    //: /sn:0 {0}(-323,371)(-393,371){1}
wire w14;    //: /sn:0 {0}(271,76)(271,161)(394,161)(394,309){1}
wire w4;    //: /sn:0 {0}(529,366)(451,366){1}
wire w15;    //: /sn:0 {0}(-427,324)(-427,273)(-167,273)(-167,328)(-125,328){1}
wire w38;    //: /sn:0 {0}(-423,15)(-423,184)(-100,184)(-100,293){1}
wire w0;    //: /sn:0 {0}(-125,369)(-166,369)(-166,362)(-209,362){1}
wire w20;    //: /sn:0 {0}(-2,293)(-2,254)(298,254)(298,340)(334,340){1}
wire w23;    //: /sn:0 {0}(345,76)(345,149)(491,149)(491,224)(561,224)(561,332){1}
wire w41;    //: /sn:0 {0}(-494,15)(-494,214)(-301,214)(-301,307){1}
wire w18;    //: /sn:0 {0}(-323,341)(-374,341)(-374,255)(-551,255)(-551,360)(-573,360){1}
wire w8;    //: /sn:0 {0}(627,109)(627,332){1}
wire w35;    //: /sn:0 {0}(-2,44)(-2,206)(362,206)(362,309){1}
wire w17;    //: /sn:0 {0}(197,294)(197,135)(200,135)(200,76){1}
wire w2;    //: /sn:0 {0}(477,109)(477,121)(452,121)(452,190)(224,190)(224,294){1}
wire w44;    //: /sn:0 {0}(-475,324)(-475,233)(-573,233)(-573,15){1}
wire w12;    //: /sn:0 {0}(110,374)(77,374)(77,358)(29,358){1}
wire w10;    //: /sn:0 {0}(-573,365)(-508,365){1}
wire w13;    //: /sn:0 {0}(110,329)(78,329)(78,238)(-235,238)(-235,307){1}
wire w5;    //: /sn:0 {0}(556,109)(556,180)(520,180)(520,273)(425,273)(425,309){1}
wire w29;    //: /sn:0 {0}(-147,44)(-147,158)(-68,158)(-68,293){1}
wire w47;    //: /sn:0 {0}(-349,15)(-349,170)(133,170)(133,294){1}
wire w26;    //: /sn:0 {0}(-76,44)(-76,134)(164,134)(164,294){1}
//: enddecls

  _GGAND2 #(6) g4 (.I0(B0), .I1(A1), .Z(w8));   //: @(627,99) /sn:0 /R:3 /anc:1 /w:[ 13 11 0 ]
  _GGAND2 #(6) g8 (.I0(B1), .I1(A0), .Z(w23));   //: @(345,66) /sn:0 /R:3 /w:[ 11 13 0 ]
  //: comment g61 @(9,29) /sn:0
  //: /line:"A0B2"
  //: /end
  //: OUT g86 (S7) @(-611,456) /sn:0 /R:3 /w:[ 1 ]
  _GGAND2 #(6) g3 (.I0(B0), .I1(A2), .Z(w5));   //: @(556,99) /sn:0 /R:3 /anc:1 /w:[ 15 11 0 ]
  _GGAND2 #(6) g13 (.I0(B2), .I1(A0), .Z(w35));   //: @(-2,34) /sn:0 /R:3 /w:[ 11 15 0 ]
  //: comment g34 @(568,89) /sn:0
  //: /line:"A2B0"
  //: /end
  //: joint g37 (A0) @(343, -207) /w:[ 6 -1 5 12 ]
  //: joint g51 (A2) @(-149, -140) /w:[ 4 -1 3 14 ]
  //: joint g55 (B2) @(-144, -17) /w:[ 4 -1 3 14 ]
  //: joint g58 (A1) @(-425, -175) /w:[ 2 -1 1 16 ]
  _GGAND2 #(6) g2 (.I0(B0), .I1(A3), .Z(w2));   //: @(477,99) /sn:0 /R:3 /anc:1 /w:[ 17 9 0 ]
  //: joint g65 (B3) @(-346, -46) /w:[ 8 -1 7 10 ]
  //: OUT g76 (S2) @(391,459) /sn:0 /R:3 /w:[ 1 ]
  FA4a g77 (.D(w2), .C(w17), .B(w26), .A(w47), .Cin(w7), .C2(w13), .C1(w12), .S0(S3));   //: @(111, 295) /sz:(136, 111) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>1 Ri0>1 Lo0<0 Lo1<0 Bo0<0 ]
  //: joint g59 (A2) @(-496, -140) /w:[ 2 -1 1 16 ]
  _GGAND2 #(6) g1 (.I0(B1), .I1(A1), .Z(w14));   //: @(271,66) /sn:0 /R:3 /w:[ 13 13 0 ]
  //: comment g72 @(-562,-1) /sn:0
  //: /line:"A3B3"
  //: /end
  //: comment g64 @(-215,25) /sn:0
  //: /line:"A3B2"
  //: /end
  _GGAND2 #(6) g11 (.I0(B2), .I1(A2), .Z(w29));   //: @(-147,34) /sn:0 /R:3 /w:[ 15 15 0 ]
  _GGAND2 #(6) g16 (.I0(B3), .I1(A2), .Z(w41));   //: @(-494,5) /sn:0 /R:3 /w:[ 15 17 0 ]
  _GGAND2 #(6) g10 (.I0(B2), .I1(A1), .Z(w26));   //: @(-76,34) /sn:0 /R:3 /w:[ 13 15 0 ]
  //: joint g28 (B0) @(480, 49) /w:[ 2 -1 1 16 ]
  //: joint g50 (A1) @(-78, -175) /w:[ 4 -1 3 14 ]
  //: OUT g78 (S3) @(178,459) /sn:0 /R:3 /w:[ 1 ]
  //: IN g19 (B3) @(-619,-46) /sn:0 /w:[ 0 ]
  //: joint g27 (B0) @(559, 49) /w:[ 4 -1 3 14 ]
  //: comment g32 @(713,90) /sn:0
  //: /line:"A0B0"
  //: /end
  _GGAND2 #(6) g6 (.I0(B1), .I1(A2), .Z(w17));   //: @(200,66) /sn:0 /R:3 /w:[ 15 13 1 ]
  //: joint g38 (A1) @(269, -175) /w:[ 6 -1 5 12 ]
  //: comment g69 @(-337,-1) /sn:0
  //: /line:"A0B3"
  //: /end
  _GGAND2 #(6) g7 (.I0(B1), .I1(A3), .Z(w6));   //: @(121,66) /sn:0 /R:3 /w:[ 17 11 0 ]
  //: IN g9 (B1) @(82,15) /sn:0 /w:[ 0 ]
  //: joint g53 (B2) @(1, -17) /w:[ 8 -1 7 10 ]
  //: joint g57 (A0) @(-351, -207) /w:[ 2 -1 1 16 ]
  FA3alt g75 (.C(w5), .B(w14), .A(w35), .Cin(w4), .C2(w20), .C1(w7), .S(S2));   //: @(335, 310) /sz:(115, 95) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ri0>1 Lo0<1 Lo1<0 Bo0<0 ]
  _GGAND2 #(6) g15 (.I0(B3), .I1(A1), .Z(w38));   //: @(-423,5) /sn:0 /R:3 /w:[ 13 17 0 ]
  //: joint g20 (B0) @(704, 49) /anc:1 /w:[ 8 -1 7 10 ]
  //: joint g31 (A3) @(475, -99) /w:[ 6 -1 5 8 ]
  //: comment g71 @(-482,-1) /sn:0
  //: /line:"A2B3"
  //: /end
  //: joint g39 (A2) @(198, -140) /w:[ 6 -1 5 12 ]
  //: joint g67 (B3) @(-491, -46) /w:[ 4 -1 3 14 ]
  //: joint g68 (B3) @(-570, -46) /w:[ 2 -1 1 16 ]
  //: comment g43 @(211,59) /sn:0
  //: /line:"A2B1"
  //: /end
  //: joint g48 (B1) @(348, 15) /w:[ 8 -1 7 10 ]
  _GGAND2 #(6) g17 (.I0(B3), .I1(A3), .Z(w44));   //: @(-573,5) /sn:0 /R:3 /w:[ 17 17 1 ]
  //: joint g25 (A0) @(699, -207) /w:[ 8 -1 7 10 ]
  //: joint g29 (A1) @(625, -175) /w:[ 8 -1 7 10 ]
  //: comment g62 @(-65,26) /sn:0
  //: /line:"A1B2"
  //: /end
  FAdD g73 (.in2(w8), .in1(w23), .CoutFAd(w4), .S(S1));   //: @(530, 333) /sz:(128, 69) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: comment g42 @(282,59) /sn:0
  //: /line:"A1B1"
  //: /end
  //: joint g52 (A3) @(-228, -99) /w:[ 2 -1 12 1 ]
  //: comment g63 @(-137,26) /sn:0
  //: /line:"A2B2"
  //: /end
  FAb g83 (.B(w15), .A(w44), .Cin(w16), .Cout(w10), .S(S6));   //: @(-507, 325) /sz:(113, 82) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  //: OUT g74 (S1) @(600,459) /sn:0 /R:3 /w:[ 1 ]
  _GGAND2 #(6) g5 (.I0(B0), .I1(A0), .Z(S0));   //: @(701,99) /sn:0 /R:3 /anc:1 /w:[ 11 11 0 ]
  //: IN g14 (B2) @(-265,-17) /sn:0 /w:[ 0 ]
  //: joint g56 (B2) @(-223, -17) /w:[ 2 -1 1 16 ]
  //: comment g44 @(132,59) /sn:0
  //: /line:"A3B1"
  //: /end
  //: joint g47 (B1) @(274, 15) /w:[ 6 -1 5 12 ]
  FA4b g79 (.D(w20), .C(w6), .B(w29), .A(w38), .Cin(w12), .C2(w15), .C1(w0), .S0(S4));   //: @(-124, 294) /sz:(152, 113) /sn:0 /p:[ Ti0>0 Ti1>1 Ti2>1 Ti3>1 Ri0>1 Lo0<1 Lo1<0 Bo0<0 ]
  //: OUT g80 (S4) @(-49,457) /sn:0 /R:3 /w:[ 1 ]
  _GGOR2 #(6) g85 (.I0(w10), .I1(w18), .Z(S7));   //: @(-584,362) /sn:0 /R:2 /w:[ 0 1 0 ]
  //: OUT g84 (S6) @(-452,456) /sn:0 /R:3 /w:[ 1 ]
  //: IN g21 (A0) @(-621,-207) /sn:0 /anc:1 /w:[ 0 ]
  //: IN g24 (A3) @(-621,-99) /sn:0 /anc:1 /w:[ 15 ]
  //: OUT g36 (S0) @(701,459) /sn:0 /R:3 /w:[ 1 ]
  //: IN g23 (A2) @(-621,-140) /sn:0 /anc:1 /w:[ 0 ]
  //: comment g41 @(356,60) /sn:0
  //: /line:"A0B1"
  //: /end
  //: joint g40 (A3) @(119, -99) /w:[ 4 -1 3 10 ]
  //: joint g54 (B2) @(-73, -17) /w:[ 6 -1 5 12 ]
  //: joint g60 (A3) @(-575, -99) /w:[ 13 -1 14 16 ]
  FA3b g81 (.C(w13), .B(w32), .A(w41), .Cin(w0), .C2(w18), .C1(w16), .S(S5));   //: @(-322, 308) /sz:(112, 98) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ri0>1 Lo0<0 Lo1<0 Bo0<0 ]
  //: IN g0 (B0) @(437,49) /sn:0 /anc:1 /w:[ 0 ]
  //: IN g22 (A1) @(-622,-175) /sn:0 /anc:1 /w:[ 0 ]
  //: joint g26 (B0) @(630, 49) /w:[ 6 -1 5 12 ]
  //: comment g35 @(487,89) /sn:0
  //: /line:"A3B0"
  //: /end
  //: joint g45 (B1) @(124, 15) /w:[ 2 -1 1 16 ]
  //: joint g46 (B1) @(203, 15) /w:[ 4 -1 3 14 ]
  //: comment g70 @(-411,-2) /sn:0
  //: /line:"A1B3"
  //: /end
  //: OUT g82 (S5) @(-265,456) /sn:0 /R:3 /w:[ 1 ]
  //: joint g66 (B3) @(-420, -46) /w:[ 6 -1 5 12 ]
  _GGAND2 #(6) g12 (.I0(B2), .I1(A3), .Z(w32));   //: @(-226,34) /sn:0 /R:3 /w:[ 17 0 0 ]
  _GGAND2 #(6) g18 (.I0(B3), .I1(A0), .Z(w47));   //: @(-349,5) /sn:0 /R:3 /w:[ 11 17 0 ]
  //: joint g30 (A2) @(554, -140) /w:[ 8 -1 7 10 ]
  //: comment g33 @(639,90) /sn:0
  //: /line:"A1B0"
  //: /end
  //: joint g49 (A0) @(-4, -207) /w:[ 4 -1 3 14 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA4b
module FA4b(C, S0, B, A, C1, C2, D, Cin);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(651,29)(658,29)(658,115){1}
input A;    //: /sn:0 {0}(587,29)(606,29)(606,115){1}
output C2;    //: /sn:0 {0}(187,398)(282,398){1}
output S0;    //: /sn:0 {0}(746,496)(695,496)(695,457){1}
input C;    //: /sn:0 {0}(696,32)(706,32)(706,115){1}
input D;    //: /sn:0 {0}(734,347)(734,297)(755,297){1}
input Cin;    //: /sn:0 {0}(881,190)(753,190){1}
output C1;    //: /sn:0 {0}(551,495)(463,495)(463,459){1}
wire w4;    //: /sn:0 {0}(659,347)(659,268){1}
wire w0;    //: /sn:0 {0}(303,401)(395,401){1}
wire w1;    //: /sn:0 {0}(571,167)(318,167)(318,396)(303,396){1}
wire w2;    //: /sn:0 {0}(632,401)(578,401)(578,301)(498,301)(498,345){1}
wire w5;    //: /sn:0 {0}(571,218)(429,218)(429,345){1}
//: enddecls

  //: IN g4 (C) @(694,32) /sn:0 /w:[ 0 ]
  //: OUT g8 (S0) @(743,496) /sn:0 /w:[ 0 ]
  //: IN g3 (B) @(649,29) /sn:0 /w:[ 0 ]
  //: IN g2 (A) @(585,29) /sn:0 /w:[ 0 ]
  FAdB g1 (.in2(D), .in1(w4), .CoutFAd(w2), .S(S0));   //: @(633, 348) /sz:(136, 108) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<1 ]
  _GGOR2 #(6) g11 (.I0(w0), .I1(w1), .Z(C2));   //: @(292,398) /sn:0 /R:2 /w:[ 0 1 1 ]
  //: OUT g10 (C1) @(548,495) /sn:0 /w:[ 0 ]
  //: OUT g6 (C2) @(190,398) /sn:0 /R:2 /w:[ 0 ]
  FAdC g9 (.in4(w5), .in3(w2), .CoutFAdC(w0), .S1(C1));   //: @(396, 346) /sz:(133, 112) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: IN g7 (D) @(757,297) /sn:0 /R:2 /w:[ 1 ]
  //: IN g5 (Cin) @(883,190) /sn:0 /R:2 /w:[ 0 ]
  FA3alt g0 (.C(C), .B(B), .A(A), .Cin(Cin), .C1(w5), .C2(w1), .S(w4));   //: @(572, 116) /sz:(180, 151) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ri0>1 Lo0<0 Lo1<0 Bo0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FAdC
module FAdC(in4, CoutFAdC, S1, in3);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output S1;    //: /sn:0 {0}(260,112)(370,112){1}
input in4;    //: /sn:0 {0}(134,142)(183,142){1}
//: {2}(187,142)(224,142)(224,114)(239,114){3}
//: {4}(185,144)(185,214)(239,214){5}
output CoutFAdC;    //: /sn:0 {0}(371,217)(260,217){1}
input in3;    //: /sn:0 {0}(134,85)(151,85){1}
//: {2}(155,85)(224,85)(224,109)(239,109){3}
//: {4}(153,87)(153,219)(239,219){5}
//: enddecls

  //: joint g4 (in3) @(153, 85) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g3 (.I0(in4), .I1(in3), .Z(CoutFAdC));   //: @(250,217) /sn:0 /w:[ 5 5 1 ]
  _GGXOR2 #(8) g2 (.I0(in3), .I1(in4), .Z(S1));   //: @(250,112) /sn:0 /w:[ 3 3 0 ]
  //: IN g1 (in4) @(132,142) /sn:0 /w:[ 0 ]
  //: OUT g6 (CoutFAdC) @(368,217) /sn:0 /w:[ 0 ]
  //: OUT g7 (S1) @(367,112) /sn:0 /w:[ 1 ]
  //: joint g5 (in4) @(185, 142) /w:[ 2 -1 1 4 ]
  //: IN g0 (in3) @(132,85) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA4a
module FA4a(C, S0, B, A, C1, C2, D, Cin);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(651,29)(658,29)(658,115){1}
input A;    //: /sn:0 {0}(587,29)(606,29)(606,115){1}
output C2;    //: /sn:0 {0}(185,398)(282,398){1}
output S0;    //: /sn:0 {0}(746,496)(695,496)(695,457){1}
input C;    //: /sn:0 {0}(696,32)(706,32)(706,115){1}
input D;    //: /sn:0 {0}(734,347)(734,297)(755,297){1}
input Cin;    //: /sn:0 {0}(881,190)(753,190){1}
output C1;    //: /sn:0 {0}(551,495)(463,495)(463,459){1}
wire w4;    //: /sn:0 {0}(659,347)(659,268){1}
wire w0;    //: /sn:0 {0}(303,401)(395,401){1}
wire w1;    //: /sn:0 {0}(571,167)(318,167)(318,396)(303,396){1}
wire w2;    //: /sn:0 {0}(632,401)(578,401)(578,301)(498,301)(498,345){1}
wire w5;    //: /sn:0 {0}(571,218)(429,218)(429,345){1}
//: enddecls

  //: IN g4 (C) @(694,32) /sn:0 /w:[ 0 ]
  //: OUT g8 (S0) @(743,496) /sn:0 /w:[ 0 ]
  //: IN g3 (B) @(649,29) /sn:0 /w:[ 0 ]
  //: IN g2 (A) @(585,29) /sn:0 /w:[ 0 ]
  FAdB g1 (.in2(D), .in1(w4), .CoutFAd(w2), .S(S0));   //: @(633, 348) /sz:(136, 108) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<1 ]
  _GGOR2 #(6) g11 (.I0(w0), .I1(w1), .Z(C2));   //: @(292,398) /sn:0 /R:2 /w:[ 0 1 1 ]
  //: OUT g10 (C1) @(548,495) /sn:0 /w:[ 0 ]
  //: OUT g6 (C2) @(188,398) /sn:0 /R:2 /w:[ 0 ]
  FAdC g9 (.in4(w5), .in3(w2), .CoutFAdC(w0), .S1(C1));   //: @(396, 346) /sz:(133, 112) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: IN g7 (D) @(757,297) /sn:0 /R:2 /w:[ 1 ]
  //: IN g5 (Cin) @(883,190) /sn:0 /R:2 /w:[ 0 ]
  FA3alt g0 (.C(C), .B(B), .A(A), .Cin(Cin), .C1(w5), .C2(w1), .S(w4));   //: @(572, 116) /sz:(180, 151) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ri0>1 Lo0<0 Lo1<0 Bo0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA
module FA(Cout, Cin, B, A, Sin);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(156,149)(201,149){1}
//: {2}(205,149)(227,149)(227,132)(242,132){3}
//: {4}(203,151)(203,281)(242,281){5}
input A;    //: /sn:0 {0}(156,118)(175,118){1}
//: {2}(179,118)(227,118)(227,127)(242,127){3}
//: {4}(177,120)(177,286)(242,286){5}
output Cout;    //: /sn:0 {0}(430,282)(511,282){1}
output Sin;    //: /sn:0 {0}(430,166)(503,166){1}
input Cin;    //: /sn:0 {0}(156,208)(251,208){1}
//: {2}(255,208)(394,208)(394,168)(409,168){3}
//: {4}(253,210)(253,241)(337,241){5}
wire w3;    //: /sn:0 {0}(358,239)(387,239)(387,279)(409,279){1}
wire w2;    //: /sn:0 {0}(263,130)(322,130)(322,161){1}
//: {2}(324,163)(367,163)(367,163)(409,163){3}
//: {4}(322,165)(322,236)(337,236){5}
wire w5;    //: /sn:0 {0}(263,284)(336,284)(336,284)(409,284){1}
//: enddecls

  _GGNAND2 #(4) g4 (.I0(B), .I1(A), .Z(w5));   //: @(253,284) /sn:0 /anc:1 /w:[ 5 5 0 ]
  _GGNAND2 #(4) g8 (.I0(w3), .I1(w5), .Z(Cout));   //: @(420,282) /sn:0 /w:[ 1 1 0 ]
  _GGXOR2 #(8) g3 (.I0(A), .I1(B), .Z(w2));   //: @(253,130) /sn:0 /anc:1 /w:[ 3 3 0 ]
  //: OUT g13 (Cout) @(508,282) /sn:0 /w:[ 1 ]
  //: IN g2 (Cin) @(154,208) /sn:0 /anc:1 /w:[ 0 ]
  //: IN g1 (B) @(154,149) /sn:0 /anc:1 /w:[ 0 ]
  //: joint g11 (Cin) @(253, 208) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g10 (.I0(w2), .I1(Cin), .Z(Sin));   //: @(420,166) /sn:0 /w:[ 3 3 0 ]
  //: joint g6 (B) @(203, 149) /anc:1 /w:[ 2 -1 1 4 ]
  _GGNAND2 #(4) g7 (.I0(w2), .I1(Cin), .Z(w3));   //: @(348,239) /sn:0 /w:[ 5 5 0 ]
  //: joint g9 (w2) @(322, 163) /w:[ 2 1 -1 4 ]
  //: joint g5 (A) @(177, 118) /anc:1 /w:[ 2 -1 1 4 ]
  //: IN g0 (A) @(154,118) /sn:0 /anc:1 /w:[ 0 ]
  //: OUT g12 (Sin) @(500,166) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FAdB
module FAdB(in2, CoutFAd, S, in1);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(134,85)(151,85){1}
//: {2}(155,85)(224,85)(224,109)(239,109){3}
//: {4}(153,87)(153,219)(239,219){5}
input in2;    //: /sn:0 {0}(134,142)(183,142){1}
//: {2}(187,142)(224,142)(224,114)(239,114){3}
//: {4}(185,144)(185,214)(239,214){5}
output CoutFAd;    //: /sn:0 {0}(371,217)(260,217){1}
output S;    //: /sn:0 {0}(260,112)(370,112){1}
//: enddecls

  //: joint g4 (in1) @(153, 85) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g3 (.I0(in2), .I1(in1), .Z(CoutFAd));   //: @(250,217) /sn:0 /w:[ 5 5 1 ]
  _GGXOR2 #(8) g2 (.I0(in1), .I1(in2), .Z(S));   //: @(250,112) /sn:0 /w:[ 3 3 0 ]
  //: IN g1 (in2) @(132,142) /sn:0 /w:[ 0 ]
  //: OUT g6 (CoutFAd) @(368,217) /sn:0 /w:[ 0 ]
  //: OUT g7 (S) @(367,112) /sn:0 /w:[ 1 ]
  //: joint g5 (in2) @(185, 142) /w:[ 2 -1 1 4 ]
  //: IN g0 (in1) @(132,85) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

